
//Количество байтов, которые передаются по dat линиям
typedef bit [8:0] type_data4_count;